module gameFSM (reset, clock, collided, reached_screen_end, user_input, col);

    localparam S_BEGIN = 2'b00,
                S_CONTINUE = 2'b01,
                S_LOST = 2'b10,
                S_WON = 2'b11 ;

    input collided, reached_screen_end, user_input; //user input is a boolean value (=1 when user is providing some input )
    input reset, clock;
    reg [1:0] current_state, next_state;
	output reg [2:0] col;

    always @ (*)  //next state logic
    begin : state_table
        if (!reset) begin
	 next_state = S_BEGIN;
	col <= 3'b110;
        case (current_state)
            S_BEGIN : next_state = user_input ? S_CONTINUE : S_BEGIN;

            S_CONTINUE : begin
                if (collided)
                    next_state = S_LOST;
                else if (reached_screen_end)
                    next_state = S_WON;
            end

            S_LOST : begin
		next_state = S_BEGIN;
		col <= 3'b100;
		end
            S_WON : begin
		next_state = S_BEGIN;
		col <= 3'b010;
		end

            default : next_state = S_BEGIN;
        endcase
    end
	end 

//what output to give from this module?
	// State update logic
    always @ (posedge clock) begin
        if (!reset) 
            current_state <= S_BEGIN;
        else 
            current_state <= next_state;
    end
endmodule
